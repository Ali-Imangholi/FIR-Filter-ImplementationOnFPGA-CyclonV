module async_receiver(
    input clk,
    input RxD,
    output reg RxD_data_ready = 0,
    output reg [7:0] RxD_data = 0  // data received, valid only (for one clock cycle) when RxD_data_ready is asserted
);

parameter ClkFrequency = 50000000;
parameter Baud = 115200;
parameter Oversampling = 4;	// needs to be a power of 2

reg [3:0] RxD_state = 0;
wire sample;
reg [1:0] count = 0;
reg cout;

BaudTickGen #(ClkFrequency, Baud, Oversampling) tickgen(.clk(clk), .enable((RxD_state==4'b0000)), .tick(sample));
//assign RxD_data_ready = (RxD_state == 4'b1011);

always @(posedge clk)
begin

      
 

    if((RxD_state == 4'b0000) & !RxD)
        RxD_data[0]= RxD;
        
    else if((RxD_state > 4'b0010) & cout)
        RxD_data <= { RxD, RxD_data[7:1]};

	 case(RxD_state)
        4'b0000: if(!RxD) RxD_state <= 4'b0001;
        4'b0001: if(count == 2'b10) RxD_state <= 4'b0010;  // start bit
        4'b0010: if(cout) RxD_state <= 4'b0011;  // start bit sampling
        4'b0011: if(cout) RxD_state <= 4'b0100;  // bit 0
        4'b0100: if(cout) RxD_state <= 4'b0101;  // bit 1
        4'b0101: if(cout) RxD_state <= 4'b0110;  // bit 2
        4'b0110: if(cout) RxD_state <= 4'b0111;  // bit 3
        4'b0111: if(cout) RxD_state <= 4'b1000;  // bit 4
        4'b1000: if(cout) RxD_state <= 4'b1001;  // bit 5
        4'b1001: if(cout) RxD_state <= 4'b1010;  // bit 6
        4'b1010: begin if(cout) RxD_state <= 4'b1011; end // bit 7
        4'b1011: begin if(sample) RxD_state <= 4'b0000;  RxD_data_ready=1; end  // stop1
        default: if(RxD) RxD_state <= 4'b0000;
     endcase  
end

always@( sample)begin

      if (RxD_state == 4'b0000) begin
	count = 2'b00;
	cout = 0; end 
     else if ( sample)begin
      
	count = count + 1;
	cout = 0; end

     if (count == 2'b11 & sample)
	  cout = 1'b1;
	  else if(count == 2'b11 & ~sample)
     cout = 1'b0;
end


endmodule

